library ieee;
use ieee.std_logic_1164.all;

entity datapath is
    generic (N: integer := 18);
    port (
    );
end entity;

architecture operative_block of datapath is
end architecture;































